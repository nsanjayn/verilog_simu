module INV_X1 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
