module INV_X8 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
