module INV_X4 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
