module LOGIC1_X1 (Z);
  output Z;

  buf(Z, 1);
endmodule
