module XOR2_X2 (A, B, Z);
  input A;
  input B;
  output Z;

  xor(Z, A, B);


endmodule
