module FILLCELL_X16 ();

endmodule
