module ANTENNA_X1 (A);
  input A;

endmodule
