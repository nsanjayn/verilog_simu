module INV_X16 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
