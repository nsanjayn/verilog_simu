module FILLCELL_X2 ();

endmodule
