module FILLCELL_X4 ();

endmodule
