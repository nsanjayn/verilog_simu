module LOGIC0_X1 (Z);
  output Z;

  buf(Z, 0);
endmodule
