module CLKBUF_X2 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
