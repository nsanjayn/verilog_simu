module BUF_X32 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
