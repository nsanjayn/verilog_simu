module FILLCELL_X32 ();

endmodule
