module FILLCELL_X8 ();

endmodule
