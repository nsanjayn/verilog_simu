module INV_X2 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
