module BUF_X8 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
