module FILLCELL_X1 ();

endmodule
