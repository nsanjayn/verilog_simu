module BUF_X4 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
