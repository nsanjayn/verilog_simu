module BUF_X16 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
