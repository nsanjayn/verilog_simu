module INV_X32 (A, ZN);
  input A;
  output ZN;

  not(ZN, A);


endmodule
