module CLKBUF_X1 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
