module CLKBUF_X3 (A, Z);
  input A;
  output Z;

  buf(Z, A);


endmodule
